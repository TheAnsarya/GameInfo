CDLv2�%nP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    		    	       	                       		                 	                    	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            			      		                                                	                  	                       		                                                                        				                       			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  			 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                        	   	                                                                                                                             			              	                                                                                         		                                                                                                                                                                                           		                                                          		         	        	          	                                                                              	                                    	                                								   	                                                                                                                                                            	              		    						                                                                               		                                                                                                                           		                                              				      	     					   		                                                                                      	                                             		            	        	 	                                                   				     	 													              		                	                                                                                                                	  	           	             					                                                                                                                                                                                  		    		                                	                                                                   	                   		                                                                          				                                                                              				  		  		 		  						 		    		                                                                                                                						 										  					                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                                                                                                                                                                                                       		                  	                                      		                                                                                                                        	                                	                             	        	                                                                                                                                                                                                                                                                                                                                                                                                                                       				                                                                                                                                                                                       		                                                                                                                                                  	                                                                                     						  	                                                                                                                                                                      	                                                                                                                                                                                                                                                                                                                                           	                            	      	                                                                                                                                   		                                                                   	                                                                                                                                	                                               			                     	                        	          	                                                   	        	                                                                                                                                                                                                                                                                                                                                                          			                                                                        						                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                			                                                                                                                                                                                           	     		        	      				  	                                                                                                         				                                  			       	                                                                  	                                                                	                                        		                                                                                                                                                                                                                                                                                		                                                                                         	                                                                                                                        		          	                                                                       				    		                                                                               	                                			                            	                                                                            	                                     	                                                                      	   	       				  	                      	                                                                                                                                                                                                                       	                                                                                                                                                                                                                                                                               		                                                                     	                                                       	                               	    	                                                                                     				           	  	                      	                          	        	                                                                                                                                                                                                                                                                                                                                                                                                  		                                                    	                                                                                 	            	           	                                                                           	                                                              	                                                    	                                  	                                                 				                      	                                       			                                                    	                                                     			       	                 	                                                                                                                                                                                                                                                                                                                                                                                   	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                           	               	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        	                                                                                     	                                      	                                                                                                                                                                                                             					  					            		                                               	            	                                           	  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       		                                                                                                                                                                                            						                                                                                                                                					            	       	    	                                                                                                                                                                                                                                                                                          		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	                                                                                                                          	                                                                                                        	        		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	                                                                           			                                  	                            					   	    			              		                                                                                         									                                                                    			    		                            	            	                          					                                     					       		                                                    	                                                                                                                                                                                                                             					                                                               	                    	   	                                                  	              		              	                                                   				       			   							                                                               	                                                                                 			                                                               	                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                             				       	             			                        	                                                                                                                      	                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	         			                           		                     			             		    	    				               			    				           	                                    			    			                                                                       		                                                                                                                                                		                     								         	          	                        	                                                    	                                                                            	    	    	                                                                                                                                                       	                                                                                                            	                                                                                                                                                                                                                      	           		                	                                                             	                                       	                                                                                                                         	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                 	                                                                                                                                                                                                               		             				                    	                                                                                 		                        		      				       	                                  	           		                          	                             		                          	                                                                                                                                                         				                                                                                                                                                                              	          		 			                           	                                                                         			   	   	        	               	                        	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	                                                 		                                                        	        		          		 		                                                                                                                                                                                       			                                                                                              					  		  												                 					                  	             			  				                      			                    		         			 			    	    	        			                	  									  			    		      		    		  			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	                                                         		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 				                     				                        								                          			                	 	   	                                                                                     		                                                                                                                                                                                                                                                    	                                                                         	                                                                                                                                                                                                                                                                                                   		                                                                                                                                                                                                                     	   		                                                                                                                                                                                                                                                                             	 			                                         					                                                   				                                           		                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	                                                                        	                         					    	  		                                                                                               		    	                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                         	                   				                                                                                                            	     							             	                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	                                                                                                          	             	    													                                              					 	         	               	                                                                                                                                        		      	                                         				                			        			  	                             	    			                            			                                                                                                                                                                                                  	  		         		     	     		                            	                             	                                                                                                 	                   		               	   	   	   					         	  	                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                 	                                                    	                                                                                                   		                             	  	            		                                                                                                                                                              		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	 		   			     			             		  				         					                          		       				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	                       				                                                                                                                                                                                                                                                                                                             	                                                                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	             	   	      		                        		   									                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          								    											                							                   	                                                        		                                       								                                                                                                                                                                                                                                                                           	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	    		                                            	           									  		  	  							        	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                		              		    		                        		      			        	                                              	                          		                                                                                                                                                                                                                                                                                                                                                                                                                                                           	                                                                                                                                          		          	                               				                			                                    		          		                  	         				                     	     	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	     		  						                                                                                                   	  				   																		                               							 																				                  													                                                                                                                                	                  		                                               					                                                                                                                                                                                                                                                             			                                                		          	                                        		    		               			                                                                                                  	                                                                                                      	                                    		                                                                                                                                                                                         	 						  			                                                                                                             	    		                      	                              	                       				 	                        	                                                                                                                                                                                                                                                               		                          	         									              	                                   	                                                      	                                                                                                                												                                                                                                      					      						        			                   			             	                      		                                     	                        		                                        					           			         	        	       							              	        	  		  				                                                                                                                                                                                                                                                                                                                                                                                                                                                                     					          		              	                  		     					  		     		                                                                                                                     								                               	                      	                                                                                                                                                                											                                                                                                                       	                                                                           			                                                                                                                                                                                                 	                       	                                                                                                                                                    			      		                                                      	                                                                                        			  			  				                                                                                                                                                    					                                                                                                                       		                                                                                                          			   		      	         	                                                                                                                                                                  		                               			                    				                               			                                                                                                                      			  	                           	           	              		    					                                                                               		                                                                                                                           		                                              			      				       				                  	                                             		      			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          				     	 					                 		     								                		                                         		                  	  	  	           	             					                                                                                                                                                                                          	    	                                                                                                                      				                                                                                                    		                                                  	                              	                         		  			             	                                                                           		                                                                                                                                                                                           										                                                                                                                                                                                                                  		                                                            
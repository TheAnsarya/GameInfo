CDLv2�%nP                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   		    	       	                       		                  	                    	 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            			      		                                                                	                      	                       		                                                                        				                       			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  			 	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                        	   	                                                                                                                             			              	                                                                                         		                                                                                                                                                                                           		                                                          		         	        	          	                                                                              	                                    	                                								   	                                                                                                                                                            	              		    						                                                                               		                                                                                                                           		                                              				      	     					   		                                                                                      	                                             		            	        	 	                                                 	  				     	 													              		                	                                                                                                                	  	           	             					                                                                                                                                                                                  		    		                                	                                                                   	                   		                                                                          				                                                                              					  		  		 		  						 		    		                                                                                                                						 										  					                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       	                                                                                                                                                                                                                       		                  	                                      		                                                                                                                        	                                	                             	        	                      	                                                                                                                                                                                                                                                                                                                                                                                                                  				                                                                                                                                                                                       		                                                                                                                                                       	                                                                                     						  	                                                                                                                                                                      	                                                                                                                                                                                                                                                                                                                                              	                            	      	                                                                                                                                                                                 		                                                                   	                                                                                                                                 	                                               			                     	                        	          	                                                   	        	                                                                                                                                                                                                                                                                                                                                                          			                                                                        				        			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                			                                                                                                                                                                                           	     		        	      				  	                                                                                                         				                                     			       	                                                                  	                                          	                                      	                                        		                                                                                                                                                                                                                                                                                		                                                                                         	                                                                                                                        		          	                                                                       				    		                                                                               	                                			                            	                                                                            	                                          	                                                                                    	   	       				  	                      	                                                                                                                                                                                                                       	                                                                                                                                                                                                                                                                                             		                                                                     	                                                                        	                                                  	    	                                                                                     				           	  	                      	                          	        	                                                                                                                                                                                                                                                                                                                                                                                                        		                                                    	                                                                                 	            	           	                                                                           	                                                    	          	                                                    	                                  	                                                 				                      	                                       			                                                    	                                                     			             	                 	                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                           	               	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        	                                                                                     	                                      	                                                                                                                                                                                                             					  					            		                                               	            	                                           	  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       		                                                                                                                                                                                                    						                                                                                                                                					            	       	    	                                                                                                                                                                                                                                                                                           		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              	                                                                                                                             	                                                                                                        	        		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	                                                                           			                                  	                            					   	    			              		                                                                                                                                       									                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	            	                          					                                     					       		                                                    	                                                                                                                                                                                                                             					                                                               	                    	   	                                                  	              		              	                                                   				       			   							                                                               	                                                                                 			                                                               	                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                             				       	             			                        	                                                                                                                      	                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	         			                           		                     			             		    	    				               			    				           	                                    			    			                                                                       		                                                                                                                                                		                     								         	          	                        	                                                    	                                                                            	    	    	                                                                                                                                                       	                                                                                                            	                                                                                                                                                                                                                      	           		                	                                                             	                                       	                                                                                                                         	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                 	                                                                                                                                                                                                               		             				                    	                                                                                 		                        		      				       	                                  	           		                          	                             		                          	                                                                                                                                                         				                                                                                                                                                                              	          		 			                           	                                                                         			   	   	        	               	                        	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   	                                                 		                                                        	        		          		 		                                                                                                                                                                                       			                                                                                              					  		  												                 					                  	             			  				                      			                    		         			 			    	    	        			                	  										  				    		      		    		  			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	                                                         		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             				                     				                        								                          			                	 	   	                                                                                     		                                                                                                                                                                                                                                                    	                                                                         	                                                                                                                                                                                                                                                                                                   		                                                                                                                                                                                                                     	   		                                                                                                                                                                                                                                                                             	 			                                         					                                                   				                                           		                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	                                                                        	                         					    	  		                                                                                               		    	                                                                                                                                                                                                                                                  	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	                   				                                                                                                                      	     							             	                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         	                                                                                                          	             	    														                                              					 	         	               	                                                                                                                                        		      	                                         				                			        			  	                             	    			                            			                                                                                                                                                                                                          	  		         		     	     		                            	                             	                                                                                                 	                   		               	   	   	   					         	  	                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    	                 	                                                    	                                                                                                   		                             	  	              		                                                                                                                                                              		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     	  		   			     			             		  				         					                                                       		       				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                	                       				                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	             	   	      		                        		   									                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          								    											                							                   	                                                        		                                       								                                                                                                                                                                                                                                                                           	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	    		                                            	           									  		  	  							        	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                		              		    		                        		      			        	                                                  	                          		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           	                                                                                                                                          		          	                               				                			                                    		          		                  	         				                     	     	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	     		  						                                                                                                   	  				   																		                               							 																				                  													                                                                                                                                 	                                          		                                               					                                                                                                                                                                                                                                                             			                                                		          	                                              		             		               			                                                                                                  	                                                                                                      	                                    		                                                                                                                                                                                         	 						  			                                                                                                               	    		                      	                              	                       				 	                        	                                                                                                                                                                                                                                                               		                          	         									              	                                   	                                                      	                                                                                                                												                                                                                                      					      						        			                   			             	                      		                                     	                        		                                        					           			         	        	       							              	        	  		  				                                                                                                                                                                                                                                                                                                                                                                                                                                                                     					          		              	                  		     					  		     		                                                                                                                     								                               	                      	                                                                                                                                                                 											                                                                                                                       	                                                                           				                                                                                                                                                                                                        	                       	                                                                                                                                                                   			      		                                                      	                                                                                        			  			  				                                                                                                                                                    					                                                                                                                                     		                                                                                                          			   		      	         	                                                                                                                                                                  			                               			                    					                               			                                                                                                                      			  	                           	           	              		    					                                                                               		                                                                                                                           		                                              			      				       				                  	                                             		      			                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          				     	 					                 		     								                		                                         		                  	  	  	           	             					                                                                                                                                                                                          	    	                                                                                                                      				                                                                                                    		                                                  	                              	                         		  			             	                                                                           		                                                                                                                                                                                           										                                                                                                                                                                                                                  		                                                            